* D:\Analog_VLSI\eSIM\FOSSEE\eSim\library\SubcircuitLibrary\4_OR_subckt\4_OR_subckt.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/25/22 18:51:57

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_X1-Pad3_ NOR		
X2  Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_X2-Pad3_ NOR		
X3  Net-_X1-Pad3_ Net-_X2-Pad3_ Net-_U1-Pad5_ NAND		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ PORT		

.end
