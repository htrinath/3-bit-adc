* D:\Analog_VLSI\eSIM\FOSSEE\eSim\library\SubcircuitLibrary\comparator_subckt\comparator_subckt.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/24/22 14:24:04

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M6  Net-_M3-Pad2_ Net-_M1-Pad2_ Net-_M3-Pad1_ Net-_M3-Pad2_ eSim_MOS_P		
M3  Net-_M3-Pad1_ Net-_M3-Pad2_ Net-_M1-Pad1_ Net-_M3-Pad2_ eSim_MOS_P		
M9  Net-_M3-Pad1_ Net-_M9-Pad2_ Net-_M10-Pad1_ Net-_M3-Pad2_ eSim_MOS_P		
M8  Net-_M10-Pad1_ Net-_M2-Pad1_ Net-_M11-Pad1_ Net-_M3-Pad2_ eSim_MOS_P		
M4  Net-_M1-Pad1_ Net-_M11-Pad1_ Net-_M2-Pad1_ Net-_M3-Pad2_ eSim_MOS_P		
M7  Net-_M11-Pad1_ Net-_M2-Pad1_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
M5  Net-_M2-Pad1_ Net-_M11-Pad1_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
M2  Net-_M2-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
M10  Net-_M10-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
M11  Net-_M11-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
M13  Net-_M13-Pad1_ Net-_M11-Pad1_ Net-_M12-Pad1_ Net-_M13-Pad1_ eSim_MOS_P		
M12  Net-_M12-Pad1_ Net-_M11-Pad1_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
U1  Net-_M3-Pad2_ Net-_M9-Pad2_ Net-_M1-Pad2_ Net-_M13-Pad1_ Net-_M1-Pad3_ Net-_M12-Pad1_ PORT		

.end
