* D:\Analog_VLSI\eSIM\FOSSEE\eSim\library\SubcircuitLibrary\4x2_priority_encoder_subckt\4x2_priority_encoder_subckt.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/28/22 21:02:39

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X2  Net-_X1-Pad2_ Net-_U1-Pad3_ Net-_X2-Pad3_ AND		
X3  Net-_X2-Pad3_ Net-_U1-Pad1_ Net-_U1-Pad1_ Net-_U1-Pad6_ OR		
X1  Net-_U1-Pad2_ Net-_X1-Pad2_ inverter		
X4  Net-_U1-Pad1_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad5_ OR		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ ? Net-_U1-Pad5_ Net-_U1-Pad6_ PORT		

.end
