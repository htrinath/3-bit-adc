* D:\Analog_VLSI\eSIM\FOSSEE\eSim\library\SubcircuitLibrary\NAND_subckt\NAND_subckt.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/25/22 13:57:44

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad1_ eSim_MOS_P		
M4  Net-_M1-Pad1_ Net-_M3-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad1_ eSim_MOS_P		
M2  Net-_M1-Pad3_ Net-_M1-Pad2_ Net-_M2-Pad3_ Net-_M2-Pad3_ eSim_MOS_N		
M3  Net-_M2-Pad3_ Net-_M3-Pad2_ GND GND eSim_MOS_N		
v1  Net-_M1-Pad1_ GND DC		
U1  Net-_M1-Pad2_ Net-_M3-Pad2_ Net-_M1-Pad3_ PORT		

.end
