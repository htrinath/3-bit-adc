* D:\Analog_VLSI\eSIM\FOSSEE\eSim\library\SubcircuitLibrary\buffer_subckt\buffer_subckt.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/24/22 16:41:07

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M2  Net-_M2-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad1_ Net-_M2-Pad1_ eSim_MOS_P		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
M4  Net-_M2-Pad1_ Net-_M1-Pad1_ Net-_M3-Pad1_ Net-_M2-Pad1_ eSim_MOS_P		
M3  Net-_M3-Pad1_ Net-_M1-Pad1_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
U1  Net-_M1-Pad2_ Net-_M2-Pad1_ Net-_M1-Pad3_ Net-_M3-Pad1_ PORT		

.end
